module processor();


endmodule 